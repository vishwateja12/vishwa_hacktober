magic
tech scmos
timestamp 1619167648
<< nwell >>
rect -18 -7 30 26
<< ntransistor >>
rect -7 -33 -5 -23
rect 15 -33 17 -23
<< ptransistor >>
rect -7 0 -5 20
rect 15 0 17 20
<< ndiffusion >>
rect -8 -33 -7 -23
rect -5 -33 -4 -23
rect 14 -33 15 -23
rect 17 -33 18 -23
<< pdiffusion >>
rect -8 0 -7 20
rect -5 0 -4 20
rect 14 0 15 20
rect 17 0 18 20
<< ndcontact >>
rect -12 -33 -8 -23
rect -4 -33 0 -23
rect 10 -33 14 -23
rect 18 -33 22 -23
<< pdcontact >>
rect -12 0 -8 20
rect -4 0 0 20
rect 10 0 14 20
rect 18 0 22 20
<< polysilicon >>
rect -7 20 -5 23
rect 15 20 17 23
rect -7 -23 -5 0
rect 15 -23 17 0
rect -7 -37 -5 -33
rect 15 -37 17 -33
<< polycontact >>
rect -11 -13 -7 -9
rect 11 -20 15 -16
<< metal1 >>
rect -18 47 30 50
rect -12 20 -8 47
rect 10 20 14 47
rect -18 -13 -11 -9
rect -18 -20 11 -16
rect 10 -58 14 -33
rect -18 -61 30 -58
<< metal2 >>
rect -4 -10 0 20
rect 18 -10 22 20
rect -4 -13 30 -10
rect -12 -40 -8 -23
rect -4 -33 0 -13
rect 18 -40 22 -23
rect -12 -43 22 -40
<< labels >>
rlabel metal1 -18 47 30 50 5 vdd
rlabel metal1 -18 -61 30 -58 1 gnd
rlabel metal1 -18 -13 -7 -9 1 A
rlabel metal1 -18 -20 15 -16 1 B
rlabel metal2 -4 -13 30 -10 1 Y
rlabel metal2 -4 -23 0 -13 1 Y
rlabel metal2 18 -10 22 0 1 Y
rlabel metal2 -4 -10 0 0 1 Y
rlabel metal2 -12 -43 22 -40 1 Z
rlabel metal2 -12 -43 -8 -33 1 Z
rlabel metal2 18 -43 22 -33 1 Z
<< end >>
