magic
tech scmos
timestamp 1618809773
<< nwell >>
rect -22 -3 50 30
<< ntransistor >>
rect -9 -30 -7 -20
rect 14 -30 16 -20
rect 35 -30 37 -20
<< ptransistor >>
rect -9 3 -7 23
rect 14 3 16 23
rect 35 3 37 23
<< ndiffusion >>
rect -10 -30 -9 -20
rect -7 -30 -6 -20
rect 13 -30 14 -20
rect 16 -30 17 -20
rect 34 -30 35 -20
rect 37 -30 38 -20
<< pdiffusion >>
rect -10 3 -9 23
rect -7 3 -6 23
rect 13 3 14 23
rect 16 3 17 23
rect 34 3 35 23
rect 37 3 38 23
<< ndcontact >>
rect -14 -30 -10 -20
rect -6 -30 -2 -20
rect 9 -30 13 -20
rect 17 -30 21 -20
rect 30 -30 34 -20
rect 38 -30 42 -20
<< pdcontact >>
rect -14 3 -10 23
rect -6 3 -2 23
rect 9 3 13 23
rect 17 3 21 23
rect 30 3 34 23
rect 38 3 42 23
<< polysilicon >>
rect -9 23 -7 26
rect 14 23 16 26
rect 35 23 37 26
rect -9 -20 -7 3
rect 14 -20 16 3
rect 35 -20 37 3
rect -9 -37 -7 -30
rect 14 -37 16 -30
rect 35 -37 37 -30
<< polycontact >>
rect -13 -9 -9 -5
rect 10 -16 14 -12
rect 31 -12 35 -8
<< metal1 >>
rect -22 46 50 49
rect 9 23 13 46
rect 30 23 34 46
rect -27 -9 -13 -5
rect 38 -8 42 3
rect 27 -12 31 -8
rect 38 -12 56 -8
rect -27 -16 10 -12
rect 38 -20 42 -12
rect -14 -59 -10 -30
rect 9 -59 13 -30
rect 30 -59 34 -30
rect -22 -62 50 -59
<< m2contact >>
rect 22 -12 27 -7
<< metal2 >>
rect -14 27 21 30
rect -14 3 -11 27
rect -6 -9 -2 23
rect 17 3 21 27
rect -6 -12 22 -9
rect -6 -30 -3 -12
rect 17 -30 20 -12
<< labels >>
rlabel metal1 -22 -62 50 -59 1 gnd
rlabel metal1 -27 -9 -9 -5 1 A
rlabel metal1 -27 -16 14 -12 1 B
rlabel metal2 -6 -12 22 -9 1 Y_bar
rlabel metal1 27 -12 35 -8 1 Y_bar
rlabel metal1 42 -12 56 -8 1 Y
rlabel metal2 -14 27 21 30 1 Z
rlabel metal1 -22 46 50 49 5 vdd
<< end >>
