* SPICE3 file created from nand.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale=0.09u
.global vdd gnd

Vdd vdd gnd 'SUPPLY'

Vin_a A gnd pulse 0 1.8 0 100ps 100ps 5ns 10ns
Vin_b B gnd pulse 0 1.8 0 100ps 100ps 10ns 20ns

M1000 Y A vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1001 Z B gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1002 Y A Z Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1003 Y B vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0

.tran 0.1n 100n

.control

set hcopypscolor = 1
set color0 = white
set color1 = black

run

plot v(A)
plot v(B)
plot v(Y)
.endc

