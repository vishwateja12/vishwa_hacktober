magic
tech scmos
timestamp 1632562973
<< nwell >>
rect -31 2 -5 19
rect 1 2 65 20
rect 92 -34 144 -18
rect -45 -79 -12 -61
rect -26 -143 0 -126
rect 6 -143 70 -125
rect 97 -179 149 -163
rect -40 -224 -7 -206
rect -23 -288 3 -271
rect 9 -288 73 -270
rect 100 -324 152 -308
rect -37 -369 -4 -351
rect -15 -426 11 -409
rect 17 -426 81 -408
rect 108 -462 160 -446
rect -29 -507 4 -489
<< ntransistor >>
rect -19 -12 -17 -8
rect 14 -34 16 -30
rect 29 -34 31 -30
rect 39 -34 41 -30
rect 50 -34 52 -30
rect -32 -93 -30 -89
rect 103 -56 105 -52
rect 113 -56 115 -52
rect 131 -56 133 -52
rect -14 -157 -12 -153
rect 19 -179 21 -175
rect 34 -179 36 -175
rect 44 -179 46 -175
rect 55 -179 57 -175
rect -27 -238 -25 -234
rect 108 -201 110 -197
rect 118 -201 120 -197
rect 136 -201 138 -197
rect -11 -302 -9 -298
rect 22 -324 24 -320
rect 37 -324 39 -320
rect 47 -324 49 -320
rect 58 -324 60 -320
rect -24 -383 -22 -379
rect 111 -346 113 -342
rect 121 -346 123 -342
rect 139 -346 141 -342
rect -3 -440 -1 -436
rect 30 -462 32 -458
rect 45 -462 47 -458
rect 55 -462 57 -458
rect 66 -462 68 -458
rect -16 -521 -14 -517
rect 119 -484 121 -480
rect 129 -484 131 -480
rect 147 -484 149 -480
<< ptransistor >>
rect -19 8 -17 13
rect 14 8 16 14
rect 29 8 31 14
rect 39 8 41 14
rect 50 8 52 14
rect 103 -28 105 -24
rect 113 -28 115 -24
rect 131 -28 133 -24
rect -32 -73 -30 -67
rect -14 -137 -12 -132
rect 19 -137 21 -131
rect 34 -137 36 -131
rect 44 -137 46 -131
rect 55 -137 57 -131
rect 108 -173 110 -169
rect 118 -173 120 -169
rect 136 -173 138 -169
rect -27 -218 -25 -212
rect -11 -282 -9 -277
rect 22 -282 24 -276
rect 37 -282 39 -276
rect 47 -282 49 -276
rect 58 -282 60 -276
rect 111 -318 113 -314
rect 121 -318 123 -314
rect 139 -318 141 -314
rect -24 -363 -22 -357
rect -3 -420 -1 -415
rect 30 -420 32 -414
rect 45 -420 47 -414
rect 55 -420 57 -414
rect 66 -420 68 -414
rect 119 -456 121 -452
rect 129 -456 131 -452
rect 147 -456 149 -452
rect -16 -501 -14 -495
<< ndiffusion >>
rect -22 -12 -19 -8
rect -17 -12 -16 -8
rect 12 -34 14 -30
rect 16 -34 17 -30
rect 21 -34 29 -30
rect 31 -34 32 -30
rect 36 -34 39 -30
rect 41 -34 43 -30
rect 47 -34 50 -30
rect 52 -34 53 -30
rect -34 -93 -32 -89
rect -30 -93 -29 -89
rect 102 -56 103 -52
rect 105 -56 113 -52
rect 115 -56 118 -52
rect 130 -56 131 -52
rect 133 -56 134 -52
rect -17 -157 -14 -153
rect -12 -157 -11 -153
rect 17 -179 19 -175
rect 21 -179 22 -175
rect 26 -179 34 -175
rect 36 -179 37 -175
rect 41 -179 44 -175
rect 46 -179 48 -175
rect 52 -179 55 -175
rect 57 -179 58 -175
rect -29 -238 -27 -234
rect -25 -238 -24 -234
rect 107 -201 108 -197
rect 110 -201 118 -197
rect 120 -201 123 -197
rect 135 -201 136 -197
rect 138 -201 139 -197
rect -14 -302 -11 -298
rect -9 -302 -8 -298
rect 20 -324 22 -320
rect 24 -324 25 -320
rect 29 -324 37 -320
rect 39 -324 40 -320
rect 44 -324 47 -320
rect 49 -324 51 -320
rect 55 -324 58 -320
rect 60 -324 61 -320
rect -26 -383 -24 -379
rect -22 -383 -21 -379
rect 110 -346 111 -342
rect 113 -346 121 -342
rect 123 -346 126 -342
rect 138 -346 139 -342
rect 141 -346 142 -342
rect -6 -440 -3 -436
rect -1 -440 0 -436
rect 28 -462 30 -458
rect 32 -462 33 -458
rect 37 -462 45 -458
rect 47 -462 48 -458
rect 52 -462 55 -458
rect 57 -462 59 -458
rect 63 -462 66 -458
rect 68 -462 69 -458
rect -18 -521 -16 -517
rect -14 -521 -13 -517
rect 118 -484 119 -480
rect 121 -484 129 -480
rect 131 -484 134 -480
rect 146 -484 147 -480
rect 149 -484 150 -480
<< pdiffusion >>
rect -20 8 -19 13
rect -17 8 -16 13
rect 13 8 14 14
rect 16 8 29 14
rect 31 8 32 14
rect 37 8 39 14
rect 41 8 50 14
rect 52 8 53 14
rect 102 -28 103 -24
rect 105 -28 108 -24
rect 112 -28 113 -24
rect 115 -28 118 -24
rect 122 -28 131 -24
rect 133 -28 134 -24
rect -33 -73 -32 -67
rect -30 -73 -29 -67
rect -15 -137 -14 -132
rect -12 -137 -11 -132
rect 18 -137 19 -131
rect 21 -137 34 -131
rect 36 -137 37 -131
rect 42 -137 44 -131
rect 46 -137 55 -131
rect 57 -137 58 -131
rect 107 -173 108 -169
rect 110 -173 113 -169
rect 117 -173 118 -169
rect 120 -173 123 -169
rect 127 -173 136 -169
rect 138 -173 139 -169
rect -28 -218 -27 -212
rect -25 -218 -24 -212
rect -12 -282 -11 -277
rect -9 -282 -8 -277
rect 21 -282 22 -276
rect 24 -282 37 -276
rect 39 -282 40 -276
rect 45 -282 47 -276
rect 49 -282 58 -276
rect 60 -282 61 -276
rect 110 -318 111 -314
rect 113 -318 116 -314
rect 120 -318 121 -314
rect 123 -318 126 -314
rect 130 -318 139 -314
rect 141 -318 142 -314
rect -25 -363 -24 -357
rect -22 -363 -21 -357
rect -4 -420 -3 -415
rect -1 -420 0 -415
rect 29 -420 30 -414
rect 32 -420 45 -414
rect 47 -420 48 -414
rect 53 -420 55 -414
rect 57 -420 66 -414
rect 68 -420 69 -414
rect 118 -456 119 -452
rect 121 -456 124 -452
rect 128 -456 129 -452
rect 131 -456 134 -452
rect 138 -456 147 -452
rect 149 -456 150 -452
rect -17 -501 -16 -495
rect -14 -501 -13 -495
<< ndcontact >>
rect -27 -12 -22 -8
rect -16 -12 -11 -8
rect 8 -34 12 -30
rect 17 -34 21 -30
rect 32 -34 36 -30
rect 43 -34 47 -30
rect 53 -34 57 -30
rect -38 -93 -34 -89
rect -29 -93 -25 -89
rect 98 -56 102 -52
rect 118 -56 122 -52
rect 126 -56 130 -52
rect 134 -56 138 -52
rect -22 -157 -17 -153
rect -11 -157 -6 -153
rect 13 -179 17 -175
rect 22 -179 26 -175
rect 37 -179 41 -175
rect 48 -179 52 -175
rect 58 -179 62 -175
rect -33 -238 -29 -234
rect -24 -238 -20 -234
rect 103 -201 107 -197
rect 123 -201 127 -197
rect 131 -201 135 -197
rect 139 -201 143 -197
rect -19 -302 -14 -298
rect -8 -302 -3 -298
rect 16 -324 20 -320
rect 25 -324 29 -320
rect 40 -324 44 -320
rect 51 -324 55 -320
rect 61 -324 65 -320
rect -30 -383 -26 -379
rect -21 -383 -17 -379
rect 106 -346 110 -342
rect 126 -346 130 -342
rect 134 -346 138 -342
rect 142 -346 146 -342
rect -11 -440 -6 -436
rect 0 -440 5 -436
rect 24 -462 28 -458
rect 33 -462 37 -458
rect 48 -462 52 -458
rect 59 -462 63 -458
rect 69 -462 73 -458
rect -22 -521 -18 -517
rect -13 -521 -9 -517
rect 114 -484 118 -480
rect 134 -484 138 -480
rect 142 -484 146 -480
rect 150 -484 154 -480
<< pdcontact >>
rect -25 8 -20 13
rect -16 8 -11 13
rect 8 8 13 14
rect 32 8 37 14
rect 53 8 57 14
rect 98 -28 102 -24
rect 108 -28 112 -24
rect 118 -28 122 -24
rect 134 -28 138 -24
rect -38 -73 -33 -67
rect -29 -73 -25 -67
rect -20 -137 -15 -132
rect -11 -137 -6 -132
rect 13 -137 18 -131
rect 37 -137 42 -131
rect 58 -137 62 -131
rect 103 -173 107 -169
rect 113 -173 117 -169
rect 123 -173 127 -169
rect 139 -173 143 -169
rect -33 -218 -28 -212
rect -24 -218 -20 -212
rect -17 -282 -12 -277
rect -8 -282 -3 -277
rect 16 -282 21 -276
rect 40 -282 45 -276
rect 61 -282 65 -276
rect 106 -318 110 -314
rect 116 -318 120 -314
rect 126 -318 130 -314
rect 142 -318 146 -314
rect -30 -363 -25 -357
rect -21 -363 -17 -357
rect -9 -420 -4 -415
rect 0 -420 5 -415
rect 24 -420 29 -414
rect 48 -420 53 -414
rect 69 -420 73 -414
rect 114 -456 118 -452
rect 124 -456 128 -452
rect 134 -456 138 -452
rect 150 -456 154 -452
rect -22 -501 -17 -495
rect -13 -501 -9 -495
<< polysilicon >>
rect -19 13 -17 16
rect 14 14 16 17
rect 29 14 31 17
rect 39 14 41 17
rect 50 14 52 17
rect -19 -8 -17 8
rect -19 -15 -17 -12
rect 14 -30 16 8
rect 29 -30 31 8
rect 39 -30 41 8
rect 50 -30 52 8
rect 70 -2 148 0
rect 70 -20 72 -2
rect 103 -24 105 -21
rect 113 -24 115 -20
rect 131 -24 133 -20
rect 14 -37 16 -34
rect -32 -67 -30 -64
rect -32 -89 -30 -73
rect -32 -96 -30 -93
rect 29 -102 31 -34
rect 39 -67 41 -34
rect 50 -66 52 -34
rect 79 -109 81 -45
rect 103 -52 105 -28
rect 113 -52 115 -28
rect 131 -52 133 -28
rect 103 -59 105 -56
rect 113 -59 115 -56
rect 131 -59 133 -56
rect -14 -132 -12 -129
rect 19 -131 21 -128
rect 34 -131 36 -128
rect 44 -131 46 -128
rect 55 -131 57 -128
rect -14 -153 -12 -137
rect -14 -160 -12 -157
rect 19 -175 21 -137
rect 34 -175 36 -137
rect 44 -175 46 -137
rect 55 -175 57 -137
rect 75 -147 152 -145
rect 75 -165 77 -147
rect 108 -169 110 -166
rect 118 -169 120 -165
rect 136 -169 138 -165
rect 19 -182 21 -179
rect -27 -212 -25 -209
rect -27 -234 -25 -218
rect -27 -241 -25 -238
rect 34 -247 36 -179
rect 44 -212 46 -179
rect 55 -211 57 -179
rect 84 -254 86 -190
rect 108 -197 110 -173
rect 118 -197 120 -173
rect 136 -197 138 -173
rect 108 -204 110 -201
rect 118 -204 120 -201
rect 136 -204 138 -201
rect -11 -277 -9 -274
rect 22 -276 24 -273
rect 37 -276 39 -273
rect 47 -276 49 -273
rect 58 -276 60 -273
rect -11 -298 -9 -282
rect -11 -305 -9 -302
rect 22 -320 24 -282
rect 37 -320 39 -282
rect 47 -320 49 -282
rect 58 -320 60 -282
rect 78 -292 156 -290
rect 78 -310 80 -292
rect 111 -314 113 -311
rect 121 -314 123 -310
rect 139 -314 141 -310
rect 22 -327 24 -324
rect -24 -357 -22 -354
rect -24 -379 -22 -363
rect -24 -386 -22 -383
rect 37 -392 39 -324
rect 47 -357 49 -324
rect 58 -356 60 -324
rect 87 -399 89 -335
rect 111 -342 113 -318
rect 121 -342 123 -318
rect 139 -342 141 -318
rect 111 -349 113 -346
rect 121 -349 123 -346
rect 139 -349 141 -346
rect -3 -415 -1 -412
rect 30 -414 32 -411
rect 45 -414 47 -411
rect 55 -414 57 -411
rect 66 -414 68 -411
rect -3 -436 -1 -420
rect -3 -443 -1 -440
rect 30 -458 32 -420
rect 45 -458 47 -420
rect 55 -458 57 -420
rect 66 -458 68 -420
rect 86 -430 163 -428
rect 86 -448 88 -430
rect 119 -452 121 -449
rect 129 -452 131 -448
rect 147 -452 149 -448
rect 30 -465 32 -462
rect -16 -495 -14 -492
rect -16 -517 -14 -501
rect -16 -524 -14 -521
rect 45 -530 47 -462
rect 55 -495 57 -462
rect 66 -494 68 -462
rect 95 -537 97 -473
rect 119 -480 121 -456
rect 129 -480 131 -456
rect 147 -480 149 -456
rect 119 -487 121 -484
rect 129 -487 131 -484
rect 147 -487 149 -484
<< polycontact >>
rect -23 -4 -19 0
rect 9 -11 14 -7
rect 65 -18 70 -12
rect -36 -86 -32 -82
rect 23 -102 29 -98
rect 35 -64 39 -59
rect 46 -63 50 -59
rect 52 -41 56 -37
rect 99 -42 103 -38
rect 75 -109 79 -105
rect 81 -49 85 -45
rect 109 -49 113 -45
rect 127 -41 131 -37
rect 138 -42 142 -38
rect -18 -149 -14 -145
rect 14 -156 19 -152
rect 70 -163 75 -157
rect -31 -231 -27 -227
rect 28 -247 34 -243
rect 40 -209 44 -204
rect 51 -208 55 -204
rect 57 -186 61 -182
rect 104 -187 108 -183
rect 80 -254 84 -250
rect 86 -194 90 -190
rect 114 -194 118 -190
rect 132 -186 136 -182
rect 143 -187 147 -183
rect -15 -294 -11 -290
rect 17 -301 22 -297
rect 73 -308 78 -302
rect -28 -376 -24 -372
rect 31 -392 37 -388
rect 43 -354 47 -349
rect 54 -353 58 -349
rect 60 -331 64 -327
rect 107 -332 111 -328
rect 83 -399 87 -395
rect 89 -339 93 -335
rect 117 -339 121 -335
rect 135 -331 139 -327
rect 146 -332 150 -328
rect -7 -432 -3 -428
rect 25 -439 30 -435
rect 81 -446 86 -440
rect -20 -514 -16 -510
rect 39 -530 45 -526
rect 51 -492 55 -487
rect 62 -491 66 -487
rect 68 -469 72 -465
rect 115 -470 119 -466
rect 91 -537 95 -533
rect 97 -477 101 -473
rect 125 -477 129 -473
rect 143 -469 147 -465
rect 154 -470 158 -466
<< metal1 >>
rect -56 21 179 25
rect -56 -51 -49 21
rect -25 13 -20 21
rect 32 14 37 21
rect -16 0 -11 8
rect 8 0 13 8
rect 53 0 57 8
rect -38 -4 -23 0
rect -16 -4 -3 0
rect 8 -4 57 0
rect -38 -44 -35 -4
rect -16 -8 -11 -4
rect -7 -7 -3 -4
rect -7 -11 9 -7
rect 17 -12 21 -4
rect 92 -12 96 21
rect -27 -16 -22 -12
rect -31 -19 -2 -16
rect -8 -44 -2 -19
rect 17 -18 65 -12
rect 92 -16 144 -12
rect 17 -30 21 -18
rect 98 -24 102 -16
rect 118 -24 122 -16
rect 32 -27 57 -24
rect 32 -30 36 -27
rect 53 -30 57 -27
rect 8 -38 12 -34
rect 32 -38 36 -34
rect 8 -41 36 -38
rect 43 -44 47 -34
rect 108 -37 112 -28
rect 56 -38 94 -37
rect 56 -41 99 -38
rect 90 -42 99 -41
rect 108 -41 127 -37
rect -38 -47 -13 -44
rect -8 -47 75 -44
rect -17 -50 -13 -47
rect -56 -57 -33 -51
rect -17 -53 49 -50
rect -38 -67 -33 -57
rect 46 -59 49 -53
rect -29 -82 -25 -73
rect 35 -82 38 -64
rect -54 -86 -36 -82
rect -29 -86 38 -82
rect -54 -105 -47 -86
rect -29 -89 -25 -86
rect 70 -89 75 -47
rect 85 -49 109 -45
rect 118 -52 122 -41
rect 134 -52 138 -28
rect 142 -42 148 -38
rect 98 -59 102 -56
rect 126 -59 130 -56
rect 93 -63 145 -59
rect 93 -89 97 -63
rect 56 -90 198 -89
rect -1 -93 198 -90
rect -38 -97 -34 -93
rect -1 -97 6 -93
rect -38 -101 6 -97
rect 23 -105 29 -102
rect -54 -109 75 -105
rect -51 -124 179 -120
rect -51 -196 -44 -124
rect -20 -132 -15 -124
rect 37 -131 42 -124
rect -11 -145 -6 -137
rect 13 -145 18 -137
rect 58 -145 62 -137
rect -33 -149 -18 -145
rect -11 -149 2 -145
rect 13 -149 62 -145
rect -33 -189 -30 -149
rect -11 -153 -6 -149
rect -2 -152 2 -149
rect -2 -156 14 -152
rect 22 -157 26 -149
rect 97 -157 101 -124
rect -22 -161 -17 -157
rect -26 -164 3 -161
rect -3 -189 3 -164
rect 22 -163 70 -157
rect 97 -161 149 -157
rect 22 -175 26 -163
rect 103 -169 107 -161
rect 123 -169 127 -161
rect 37 -172 62 -169
rect 37 -175 41 -172
rect 58 -175 62 -172
rect 13 -183 17 -179
rect 37 -183 41 -179
rect 13 -186 41 -183
rect 48 -189 52 -179
rect 113 -182 117 -173
rect 61 -183 99 -182
rect 61 -186 104 -183
rect 95 -187 104 -186
rect 113 -186 132 -182
rect -33 -192 -8 -189
rect -3 -192 80 -189
rect -12 -195 -8 -192
rect -51 -202 -28 -196
rect -12 -198 54 -195
rect -33 -212 -28 -202
rect 51 -204 54 -198
rect -24 -227 -20 -218
rect 40 -227 43 -209
rect -49 -231 -31 -227
rect -24 -231 43 -227
rect -49 -250 -42 -231
rect -24 -234 -20 -231
rect 75 -234 80 -192
rect 90 -194 114 -190
rect 123 -197 127 -186
rect 139 -197 143 -173
rect 147 -187 152 -183
rect 103 -204 107 -201
rect 131 -204 135 -201
rect 98 -208 150 -204
rect 98 -234 102 -208
rect 61 -235 102 -234
rect 4 -238 198 -235
rect -33 -242 -29 -238
rect 4 -242 11 -238
rect 98 -239 198 -238
rect -33 -246 11 -242
rect 28 -250 34 -247
rect -49 -254 80 -250
rect -48 -269 179 -265
rect -48 -341 -41 -269
rect -17 -277 -12 -269
rect 40 -276 45 -269
rect -8 -290 -3 -282
rect 16 -290 21 -282
rect 61 -290 65 -282
rect -30 -294 -15 -290
rect -8 -294 5 -290
rect 16 -294 65 -290
rect -30 -334 -27 -294
rect -8 -298 -3 -294
rect 1 -297 5 -294
rect 1 -301 17 -297
rect 25 -302 29 -294
rect 100 -302 104 -269
rect -19 -306 -14 -302
rect -23 -309 6 -306
rect 0 -334 6 -309
rect 25 -308 73 -302
rect 100 -306 152 -302
rect 25 -320 29 -308
rect 106 -314 110 -306
rect 126 -314 130 -306
rect 40 -317 65 -314
rect 40 -320 44 -317
rect 61 -320 65 -317
rect 16 -328 20 -324
rect 40 -328 44 -324
rect 16 -331 44 -328
rect 51 -334 55 -324
rect 116 -327 120 -318
rect 64 -328 102 -327
rect 64 -331 107 -328
rect 98 -332 107 -331
rect 116 -331 135 -327
rect -30 -337 -5 -334
rect 0 -337 83 -334
rect -9 -340 -5 -337
rect -48 -347 -25 -341
rect -9 -343 57 -340
rect -30 -357 -25 -347
rect 54 -349 57 -343
rect -21 -372 -17 -363
rect 43 -372 46 -354
rect -46 -376 -28 -372
rect -21 -376 46 -372
rect -46 -395 -39 -376
rect -21 -379 -17 -376
rect 78 -379 83 -337
rect 93 -339 117 -335
rect 126 -342 130 -331
rect 142 -342 146 -318
rect 150 -332 156 -328
rect 106 -349 110 -346
rect 134 -349 138 -346
rect 101 -353 153 -349
rect 101 -379 105 -353
rect 64 -380 198 -379
rect 7 -383 198 -380
rect -30 -387 -26 -383
rect 7 -387 14 -383
rect -30 -391 14 -387
rect 31 -395 37 -392
rect -46 -399 83 -395
rect -40 -407 179 -403
rect -40 -479 -33 -407
rect -9 -415 -4 -407
rect 48 -414 53 -407
rect 0 -428 5 -420
rect 24 -428 29 -420
rect 69 -428 73 -420
rect -22 -432 -7 -428
rect 0 -432 13 -428
rect 24 -432 73 -428
rect -22 -472 -19 -432
rect 0 -436 5 -432
rect 9 -435 13 -432
rect 9 -439 25 -435
rect 33 -440 37 -432
rect 108 -440 112 -407
rect -11 -444 -6 -440
rect -15 -447 14 -444
rect 8 -472 14 -447
rect 33 -446 81 -440
rect 108 -444 160 -440
rect 33 -458 37 -446
rect 114 -452 118 -444
rect 134 -452 138 -444
rect 48 -455 73 -452
rect 48 -458 52 -455
rect 69 -458 73 -455
rect 24 -466 28 -462
rect 48 -466 52 -462
rect 24 -469 52 -466
rect 59 -472 63 -462
rect 124 -465 128 -456
rect 72 -466 110 -465
rect 72 -469 115 -466
rect 106 -470 115 -469
rect 124 -469 143 -465
rect -22 -475 3 -472
rect 8 -475 91 -472
rect -1 -478 3 -475
rect -40 -485 -17 -479
rect -1 -481 65 -478
rect -22 -495 -17 -485
rect 62 -487 65 -481
rect -13 -510 -9 -501
rect 51 -510 54 -492
rect -38 -514 -20 -510
rect -13 -514 54 -510
rect -38 -533 -31 -514
rect -13 -517 -9 -514
rect 86 -517 91 -475
rect 101 -477 125 -473
rect 134 -480 138 -469
rect 150 -480 154 -456
rect 158 -470 163 -466
rect 114 -487 118 -484
rect 142 -487 146 -484
rect 109 -491 161 -487
rect 109 -517 113 -491
rect 72 -518 198 -517
rect 15 -521 198 -518
rect -22 -525 -18 -521
rect 15 -525 22 -521
rect -22 -529 22 -525
rect 39 -533 45 -530
rect -38 -537 91 -533
<< m2contact >>
rect 179 21 184 26
rect 198 -93 203 -88
rect 179 -124 184 -119
rect 198 -239 203 -234
rect 179 -269 184 -264
rect 198 -383 203 -378
rect 179 -407 184 -402
rect 198 -521 203 -516
<< metal2 >>
rect 179 -119 184 21
rect 179 -264 184 -124
rect 179 -402 184 -269
rect 198 -234 203 -93
rect 198 -378 203 -239
rect 198 -516 203 -383
<< labels >>
rlabel metal1 -32 -4 -32 0 1 A0
rlabel metal1 -42 -86 -42 -82 1 B0
rlabel metal1 -10 -4 -10 0 1 A0_
rlabel metal1 -22 -86 -22 -82 1 B0_
rlabel metal1 -56 -57 -33 -51 1 vdd
rlabel pdiffusion 21 8 21 14 1 D0
rlabel pdiffusion 46 8 46 14 1 E0
rlabel metal1 92 -42 92 -37 1 A0
rlabel metal1 92 -49 92 -45 1 B0
rlabel ndiffusion 109 -56 109 -52 1 F0
rlabel metal1 145 -42 145 -38 1 G0
rlabel metal1 22 -18 22 -12 1 P0
rlabel metal1 60 -18 60 -12 1 P0
rlabel metal1 120 -41 120 -37 1 C0
rlabel metal1 -38 -101 6 -97 1 gnd
rlabel metal1 -31 -19 -2 -16 1 gnd
rlabel metal1 24 -41 24 -38 1 H0
rlabel metal1 43 -27 43 -24 1 H0
rlabel metal1 92 -16 144 -12 1 vdd
rlabel metal1 93 -63 145 -59 1 gnd
rlabel metal1 -8 -47 75 -44 1 gnd
rlabel ndiffusion 114 -201 114 -197 1 H1
rlabel metal1 150 -187 150 -183 1 G1
rlabel metal1 129 -186 129 -182 1 F1
rlabel metal1 97 -194 97 -190 1 B1
rlabel metal1 97 -187 97 -182 1 A1
rlabel metal1 29 -186 29 -183 1 E1
rlabel pdiffusion 50 -137 50 -131 1 D1
rlabel pdiffusion 27 -137 27 -131 1 C1
rlabel metal1 27 -163 27 -157 1 P1
rlabel metal1 -15 -231 -15 -227 1 B1_
rlabel metal1 -40 -231 -40 -227 1 B1
rlabel metal1 -4 -149 -4 -145 1 A1_
rlabel metal1 -27 -149 -27 -145 1 A1
rlabel metal1 98 -208 150 -204 1 gnd
rlabel metal1 -3 -192 80 -189 1 gnd
rlabel metal1 -26 -164 3 -161 1 gnd
rlabel metal1 -33 -246 11 -242 1 gnd
rlabel metal1 97 -161 149 -157 1 vdd
rlabel metal1 -51 -202 -28 -196 1 vdd
rlabel metal1 -23 -309 6 -306 1 gnd
rlabel metal1 -30 -391 14 -387 1 gnd
rlabel metal1 0 -337 83 -334 1 gnd
rlabel metal1 101 -353 153 -349 1 gnd
rlabel metal1 -48 -347 -25 -341 1 vdd
rlabel metal1 100 -306 152 -302 1 vdd
rlabel metal1 -21 -294 -21 -290 1 A2
rlabel metal1 0 -294 0 -290 1 A2_
rlabel metal1 -33 -376 -33 -372 1 B2
rlabel metal1 -17 -376 -17 -372 1 B2_
rlabel metal1 33 -308 33 -302 1 P2
rlabel pdiffusion 30 -282 30 -276 1 C2
rlabel pdiffusion 54 -282 54 -276 1 D2
rlabel metal1 31 -331 31 -328 1 E2
rlabel metal1 103 -332 103 -328 1 A2
rlabel metal1 105 -339 105 -335 1 B2
rlabel metal1 127 -331 127 -327 1 F2
rlabel ndiffusion 117 -346 117 -342 1 H2
rlabel metal1 153 -332 153 -328 1 G2
rlabel metal1 161 -470 161 -466 1 G3
rlabel metal1 139 -469 139 -465 1 F3
rlabel metal1 108 -477 108 -473 1 B3
rlabel metal1 110 -470 110 -466 1 A3
rlabel metal1 74 -446 74 -440 1 P3
rlabel metal1 40 -469 40 -466 1 E3
rlabel pdiffusion 62 -420 62 -414 1 D3
rlabel pdiffusion 38 -420 38 -414 1 C3
rlabel metal1 38 -432 38 -428 1 P3
rlabel metal1 -6 -514 -6 -510 1 B3_
rlabel metal1 -24 -514 -24 -510 1 B3
rlabel metal1 7 -432 7 -428 1 A3_
rlabel metal1 -19 -432 -19 -428 1 A3
rlabel metal1 109 -491 161 -487 1 gnd
rlabel metal1 8 -475 91 -472 1 gnd
rlabel metal1 -15 -447 14 -444 1 gnd
rlabel metal1 -22 -529 22 -525 1 gnd
rlabel metal1 108 -444 160 -440 1 vdd
rlabel metal1 -40 -485 -17 -479 1 vdd
rlabel metal1 -56 21 184 25 5 vdd
rlabel metal1 -51 -124 179 -120 1 vdd
rlabel metal1 -48 -269 179 -265 1 vdd
rlabel metal1 -40 -407 179 -403 1 vdd
<< end >>
