magic
tech scmos
timestamp 1618299895
<< nwell >>
rect -47 15 138 47
<< ntransistor >>
rect -33 -18 -31 -8
rect -2 -18 0 -8
rect 29 -18 31 -8
rect 59 -18 61 -8
rect 91 -18 93 -8
rect 125 -18 127 -8
<< ptransistor >>
rect -33 21 -31 41
rect -2 21 0 41
rect 29 21 31 41
rect 59 21 61 41
rect 91 21 93 41
rect 125 21 127 41
<< ndiffusion >>
rect -34 -18 -33 -8
rect -31 -18 -30 -8
rect -3 -18 -2 -8
rect 0 -18 1 -8
rect 28 -18 29 -8
rect 31 -18 32 -8
rect 58 -18 59 -8
rect 61 -18 62 -8
rect 90 -18 91 -8
rect 93 -18 94 -8
rect 124 -18 125 -8
rect 127 -18 128 -8
<< pdiffusion >>
rect -34 21 -33 41
rect -31 21 -30 41
rect -3 21 -2 41
rect 0 21 1 41
rect 28 21 29 41
rect 31 21 32 41
rect 58 21 59 41
rect 61 21 62 41
rect 90 21 91 41
rect 93 21 94 41
rect 124 21 125 41
rect 127 21 128 41
<< ndcontact >>
rect -38 -18 -34 -8
rect -30 -18 -26 -8
rect -7 -18 -3 -8
rect 1 -18 5 -8
rect 24 -18 28 -8
rect 32 -18 36 -8
rect 54 -18 58 -8
rect 62 -18 66 -8
rect 86 -18 90 -8
rect 94 -18 98 -8
rect 120 -18 124 -8
rect 128 -18 132 -8
<< pdcontact >>
rect -38 21 -34 41
rect -30 21 -26 41
rect -7 21 -3 41
rect 1 21 5 41
rect 24 21 28 41
rect 32 21 36 41
rect 54 21 58 41
rect 62 21 66 41
rect 86 21 90 41
rect 94 21 98 41
rect 120 21 124 41
rect 128 21 132 41
<< polysilicon >>
rect -33 41 -31 44
rect -2 41 0 44
rect 29 41 31 44
rect 59 41 61 44
rect 91 41 93 44
rect 125 41 127 44
rect -33 -8 -31 21
rect -2 -8 0 21
rect 29 -8 31 21
rect 59 -8 61 21
rect 91 -8 93 21
rect 125 -8 127 21
rect -33 -28 -31 -18
rect -2 -28 0 -18
rect 29 -28 31 -18
rect 59 -28 61 -18
rect 91 -28 93 -18
rect 125 -28 127 -18
<< polycontact >>
rect -31 7 -27 11
rect -6 7 -2 11
rect 25 7 29 11
rect 61 7 65 11
rect 87 7 91 11
rect 121 7 125 11
<< metal1 >>
rect -47 64 140 67
rect -47 53 -15 56
rect -18 11 -15 53
rect -7 41 -3 64
rect 24 41 28 64
rect 86 41 90 64
rect 120 41 124 64
rect 36 30 54 34
rect 1 11 5 21
rect 94 11 98 21
rect -27 7 -6 11
rect 1 7 25 11
rect 94 7 121 11
rect 1 -8 5 7
rect 94 -8 98 7
rect -7 -41 -3 -18
rect 54 -41 58 -18
rect 86 -41 90 -18
rect 120 -41 124 -18
rect -47 -44 140 -41
<< metal2 >>
rect -38 48 131 51
rect -38 41 -35 48
rect 128 41 131 48
rect -30 5 -26 41
rect 62 5 66 41
rect -37 1 140 5
rect -30 -18 -26 1
rect 32 -18 36 1
rect 24 -35 27 -18
rect 129 -35 132 -18
rect 24 -38 132 -35
<< metal3 >>
rect -47 58 78 61
rect 75 11 78 58
rect 61 7 91 11
rect -38 -30 -35 -8
rect 62 -30 65 -8
rect -38 -33 65 -30
<< labels >>
rlabel metal2 -37 1 140 5 1 Y
rlabel metal1 -47 -44 140 -41 1 gnd
rlabel metal1 -47 64 140 67 5 vdd
rlabel metal1 -47 53 -15 56 1 A
rlabel metal1 -31 7 -2 11 1 A
rlabel metal1 -18 11 -15 56 1 A
rlabel metal1 5 7 29 11 1 A_bar
rlabel metal3 61 7 91 11 1 B
rlabel metal3 75 7 78 61 1 B
rlabel metal3 -47 58 78 61 1 B
rlabel metal1 94 7 125 11 1 B_bar
rlabel metal1 36 30 54 34 1 m
rlabel metal2 -38 48 131 51 1 l
rlabel metal3 -38 -33 65 -30 1 o
rlabel metal2 24 -38 132 -35 1 n
rlabel metal2 -30 -18 -26 1 1 Y
rlabel metal2 -30 5 -26 41 1 Y
rlabel metal2 32 -18 36 5 1 Y
rlabel metal2 62 1 66 41 1 Y
rlabel metal3 -38 -33 -35 -8 1 o
rlabel metal3 62 -33 65 -8 1 o
rlabel metal2 24 -38 27 -18 1 n
rlabel metal2 129 -38 132 -18 1 n
rlabel metal2 128 41 131 51 1 l
rlabel metal2 -38 41 -35 51 1 l
<< end >>
