magic
tech scmos
timestamp 1617951155
<< nwell >>
rect -24 -17 6 23
<< ntransistor >>
rect -10 -38 -8 -28
<< ptransistor >>
rect -10 -9 -8 11
<< ndiffusion >>
rect -11 -38 -10 -28
rect -8 -38 -7 -28
<< pdiffusion >>
rect -11 -9 -10 11
rect -8 -9 -7 11
<< ndcontact >>
rect -15 -38 -11 -28
rect -7 -38 -3 -28
<< pdcontact >>
rect -15 -9 -11 11
rect -7 -9 -3 11
<< polysilicon >>
rect -10 11 -8 14
rect -10 -28 -8 -9
rect -10 -41 -8 -38
<< polycontact >>
rect -14 -25 -10 -21
<< metal1 >>
rect -24 18 6 23
rect -15 11 -11 18
rect -7 -21 -3 -9
rect -26 -25 -14 -21
rect -7 -25 13 -21
rect -7 -28 -3 -25
rect -15 -45 -11 -38
rect -25 -50 5 -45
<< labels >>
rlabel metal1 -24 18 6 23 5 vdd
rlabel metal1 -25 -50 5 -45 1 gnd
rlabel metal1 -7 -25 13 -21 1 out
rlabel metal1 -26 -25 -10 -21 1 in
rlabel metal1 -15 11 -11 18 1 vdd
<< end >>
