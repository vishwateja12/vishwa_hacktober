* SPICE3 file created from and.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale = 0.09u
.global vdd gnd

Vdd vdd gnd 'SUPPLY'

Vin_a1 A gnd pulse 0 1.8 0 100ps 100ps 10ns 20ns
Vin_b1 B gnd pulse 0 1.8 0 100ps 100ps 5ns 10ns

M1000 Y_bar B vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=300 ps=150
M1001 Y Y_bar vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1002 Y_bar A Z Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1003 Z B gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1004 Y_bar A vdd w_n23_1# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1005 Y Y_bar gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

.tran 0.1n 100n

.control

run

plot v(A) v(B)+2 v(Y)+4

.endc
