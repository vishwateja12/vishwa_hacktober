magic
tech scmos
timestamp 1619547887
<< metal1 >>
rect 975 1417 981 1844
rect 1263 1825 1267 1843
rect 1554 1826 1558 1843
rect 1854 1828 1858 1843
rect 1206 1813 1297 1816
rect 1489 1813 1588 1816
rect 1779 1813 1885 1816
rect 1206 1702 1297 1708
rect 1489 1702 1587 1708
rect 1779 1702 1884 1708
rect 1206 1591 1297 1597
rect 1489 1591 1587 1597
rect 1779 1591 1884 1597
rect 1206 1480 1297 1486
rect 1489 1480 1587 1486
rect 1779 1480 1884 1486
rect 975 1413 1020 1417
rect 1270 1413 1302 1417
rect 1560 1413 1592 1417
rect 1859 1412 1889 1417
rect 1206 1369 1297 1375
rect 1489 1369 1587 1375
rect 1779 1369 1884 1375
rect 920 1361 995 1364
rect 1148 1361 1252 1364
rect 1424 1360 1552 1363
rect 1709 1358 1852 1362
rect 1206 1258 1297 1264
rect 1489 1258 1588 1264
rect 1779 1258 1884 1264
rect 1093 1249 1122 1252
rect 1215 1249 1312 1252
rect 1375 1251 1413 1254
rect 1503 1251 1560 1254
rect 920 1242 1029 1245
rect 1206 1147 1297 1153
rect 1489 1147 1587 1153
rect 1779 1147 1884 1153
rect 920 1052 980 1055
rect 1206 1036 1297 1042
rect 1489 1036 1588 1042
rect 1779 1036 1885 1042
rect 920 969 1019 973
rect 1277 969 1302 973
rect 1566 969 1592 973
rect 1858 969 1889 973
rect 1206 928 1297 931
rect 1489 928 1587 931
rect 1779 928 1885 931
rect 1127 778 1299 781
rect 1118 260 1122 687
rect 1127 639 1130 778
rect 1141 770 1588 773
rect 1134 685 1137 740
rect 1134 267 1137 680
rect 1141 522 1144 770
rect 1158 763 1881 766
rect 1150 559 1153 740
rect 1150 274 1153 554
rect 1158 409 1161 763
rect 1174 756 2177 759
rect 1167 463 1170 739
rect 1167 280 1170 458
rect 1174 316 1177 756
rect 1180 335 1183 739
rect 1213 680 1228 683
rect 2043 679 2095 683
rect 2043 561 2054 565
rect 1223 554 1228 557
rect 1220 458 1227 461
rect 2043 457 2056 461
rect 2062 339 2071 343
rect 1180 332 1195 335
rect 1181 286 1184 332
rect 1181 283 1841 286
rect 1167 277 1642 280
rect 1150 273 1449 274
rect 1150 271 1444 273
rect 1134 264 1245 267
rect 2091 260 2095 679
rect 1118 257 1259 260
rect 1256 236 1259 257
rect 1453 257 2095 260
rect 1453 234 1456 257
rect 2101 252 2105 561
rect 1653 249 2105 252
rect 1653 230 1656 249
rect 2111 244 2115 457
rect 1851 241 2115 244
rect 1851 227 1854 241
rect 2120 87 2124 339
rect 2115 84 2124 87
rect 2115 81 2118 84
rect 1436 66 1463 69
rect 1655 66 1672 69
rect 1864 66 1890 69
rect 2081 66 2111 69
rect 1249 28 1253 38
rect 1468 28 1471 40
rect 1677 28 1680 37
rect 1894 28 1897 40
rect 2115 28 2118 41
rect 1436 -45 1463 -39
rect 1655 -45 1672 -39
rect 1864 -45 1889 -39
rect 2081 -45 2110 -39
rect 1436 -156 1463 -150
rect 1655 -156 1672 -150
rect 1864 -156 1889 -150
rect 2081 -156 2110 -150
rect 1436 -267 1463 -261
rect 1655 -267 1672 -261
rect 1864 -267 1889 -261
rect 2081 -267 2110 -261
rect 1436 -375 1463 -372
rect 1655 -375 1672 -372
rect 1864 -375 1889 -372
rect 2081 -375 2111 -372
rect 1368 -404 1381 -400
rect 1420 -404 1443 -400
rect 1583 -404 1602 -400
rect 1641 -404 1660 -400
rect 1800 -404 1814 -400
rect 1853 -404 1868 -400
rect 2020 -404 2036 -400
rect 2075 -404 2085 -400
<< m2contact >>
rect 1262 1819 1268 1825
rect 1553 1821 1559 1826
rect 1852 1822 1859 1828
rect 1264 1413 1270 1418
rect 1554 1413 1560 1418
rect 1854 1412 1859 1418
rect 995 1360 1000 1365
rect 1143 1360 1148 1365
rect 1252 1360 1257 1365
rect 1419 1359 1424 1364
rect 1552 1358 1557 1363
rect 1703 1357 1709 1362
rect 1852 1357 1858 1362
rect 1088 1248 1093 1253
rect 1122 1248 1127 1253
rect 1210 1248 1215 1253
rect 1312 1248 1317 1253
rect 1370 1250 1375 1255
rect 1413 1250 1418 1255
rect 1498 1250 1503 1255
rect 1560 1250 1565 1255
rect 1029 1242 1034 1247
rect 980 1051 985 1056
rect 1272 969 1277 974
rect 1561 969 1566 974
rect 1853 969 1858 974
rect 1299 778 1304 783
rect 1118 687 1123 692
rect 1588 770 1593 775
rect 1133 740 1138 745
rect 1133 680 1138 685
rect 1126 634 1131 639
rect 1881 763 1886 768
rect 1149 740 1154 745
rect 1150 554 1155 559
rect 1141 517 1146 522
rect 2177 756 2182 761
rect 1166 739 1171 744
rect 1166 458 1171 463
rect 1158 404 1163 409
rect 1180 739 1185 744
rect 1226 688 1231 693
rect 1208 680 1213 685
rect 2054 561 2059 566
rect 1218 553 1223 558
rect 1215 457 1220 462
rect 2056 457 2061 462
rect 2071 339 2076 344
rect 1173 311 1178 316
rect 1841 281 1846 286
rect 1642 275 1647 280
rect 1444 268 1449 273
rect 1245 263 1250 268
rect 2101 561 2106 566
rect 1255 231 1260 236
rect 2110 457 2115 462
rect 1452 229 1457 234
rect 2119 339 2124 344
rect 1652 225 1657 230
rect 1850 222 1855 227
rect 2114 76 2119 81
rect 1249 38 1254 43
rect 1467 40 1472 45
rect 1676 37 1681 42
rect 1893 40 1898 45
rect 2114 41 2119 46
rect 1443 -404 1448 -399
rect 1660 -404 1665 -399
rect 1868 -404 1873 -399
rect 2085 -404 2090 -399
<< metal2 >>
rect 1206 1642 1228 1645
rect 1000 1361 1143 1364
rect 1030 1254 1067 1257
rect 1030 1247 1033 1254
rect 1064 1252 1067 1254
rect 1064 1249 1088 1252
rect 1127 1249 1210 1252
rect 1206 1198 1219 1201
rect 985 1052 990 1055
rect 1216 942 1219 1198
rect 1017 939 1219 942
rect 1017 916 1020 939
rect 1225 935 1228 1642
rect 1264 1418 1268 1819
rect 1489 1642 1513 1645
rect 1257 1361 1419 1364
rect 1313 1254 1350 1257
rect 1313 1253 1317 1254
rect 1347 1251 1370 1254
rect 1418 1251 1498 1254
rect 1489 1198 1502 1201
rect 1272 974 1275 1051
rect 1498 941 1502 1198
rect 1026 932 1228 935
rect 1300 938 1502 941
rect 1026 916 1029 932
rect 1300 916 1303 938
rect 1510 934 1513 1642
rect 1554 1418 1558 1821
rect 1779 1642 1798 1645
rect 1557 1359 1703 1362
rect 1561 974 1564 1250
rect 1779 1198 1790 1201
rect 1787 942 1790 1198
rect 1309 931 1513 934
rect 1592 939 1790 942
rect 1309 916 1312 931
rect 1592 916 1595 939
rect 1795 935 1798 1642
rect 1854 1418 1858 1822
rect 2076 1642 2096 1645
rect 1853 974 1857 1357
rect 2076 1198 2088 1201
rect 2085 942 2088 1198
rect 1600 932 1798 935
rect 1887 939 2088 942
rect 1600 916 1603 932
rect 1887 914 1890 939
rect 2093 934 2096 1642
rect 1895 931 2096 934
rect 1895 914 1898 931
rect 1210 777 1213 779
rect 1134 774 1213 777
rect 1134 745 1137 774
rect 1493 770 1496 777
rect 1589 775 1592 780
rect 1150 767 1496 770
rect 1150 745 1153 767
rect 1784 763 1787 780
rect 1882 768 1885 783
rect 1167 760 1787 763
rect 1167 744 1170 760
rect 2079 756 2082 778
rect 2178 761 2181 782
rect 1180 753 2082 756
rect 1180 744 1183 753
rect 1123 689 1226 692
rect 1138 680 1208 683
rect 1131 634 1209 637
rect 2059 561 2101 565
rect 1155 554 1218 557
rect 1146 517 1218 520
rect 1171 458 1215 461
rect 2061 457 2110 461
rect 1163 404 1215 407
rect 2076 339 2119 343
rect 1174 306 1177 311
rect 1245 209 1248 263
rect 1256 222 1259 231
rect 1445 213 1448 268
rect 1453 225 1456 229
rect 1445 209 1449 213
rect 1644 209 1647 275
rect 1653 220 1656 225
rect 1841 209 1844 281
rect 1851 218 1854 222
rect 1440 85 1443 87
rect 1637 85 1640 87
rect 1837 85 1840 87
rect 2035 85 2038 87
rect 1249 82 1443 85
rect 1468 82 1640 85
rect 1677 82 1840 85
rect 1894 82 2038 85
rect 1249 43 1252 82
rect 1468 45 1471 82
rect 1677 42 1680 82
rect 1894 45 1897 82
rect 2115 46 2118 76
rect 1436 -204 1447 -201
rect 1655 -204 1664 -201
rect 1864 -204 1872 -201
rect 2081 -204 2089 -201
rect 2302 -204 2317 -201
rect 1443 -399 1447 -204
rect 1660 -399 1664 -204
rect 1868 -399 1872 -204
rect 2085 -399 2089 -204
rect 2313 -387 2317 -204
<< m3contact >>
rect 990 1051 995 1056
rect 1271 1051 1276 1056
rect 1209 634 1214 639
rect 1218 517 1223 522
rect 1215 404 1220 409
rect 1173 301 1178 306
rect 1255 217 1260 222
rect 1452 220 1457 225
rect 1652 215 1657 220
rect 1850 213 1855 218
<< metal3 >>
rect 995 1052 1271 1055
rect 1214 634 1228 637
rect 1223 517 1228 520
rect 1220 404 1228 407
rect 1178 302 1195 305
rect 1256 209 1259 217
rect 1453 209 1456 220
rect 1653 209 1656 215
rect 1851 209 1854 213
use flip  flip_1
timestamp 1619247596
transform 1 0 1065 0 1 1384
box -51 -12 142 432
use flip  flip_0
timestamp 1619247596
transform 1 0 1065 0 1 940
box -51 -12 142 432
use flip  flip_3
timestamp 1619247596
transform 1 0 1348 0 1 1384
box -51 -12 142 432
use flip  flip_2
timestamp 1619247596
transform 1 0 1348 0 1 940
box -51 -12 142 432
use flip  flip_5
timestamp 1619247596
transform 1 0 1638 0 1 1384
box -51 -12 142 432
use flip  flip_4
timestamp 1619247596
transform 1 0 1638 0 1 940
box -51 -12 142 432
use flip  flip_7
timestamp 1619247596
transform 1 0 1935 0 1 1384
box -51 -12 142 432
use flip  flip_6
timestamp 1619247596
transform 1 0 1935 0 1 940
box -51 -12 142 432
use PG  PG_0
timestamp 1618762910
transform 1 0 1040 0 1 794
box -23 -17 1142 122
use CLA  CLA_0
timestamp 1618832946
transform 1 0 1252 0 1 299
box -59 -10 810 434
use sum  sum_0
timestamp 1618423665
transform 1 0 1283 0 1 94
box -40 -7 755 115
use flip  flip_8
timestamp 1619247596
transform 1 0 1295 0 -1 57
box -51 -12 142 432
use flip  flip_9
timestamp 1619247596
transform 1 0 1514 0 -1 57
box -51 -12 142 432
use flip  flip_10
timestamp 1619247596
transform 1 0 1723 0 -1 57
box -51 -12 142 432
use flip  flip_11
timestamp 1619247596
transform 1 0 1940 0 -1 57
box -51 -12 142 432
use flip  flip_12
timestamp 1619247596
transform 1 0 2161 0 -1 57
box -51 -12 142 432
use Inv  Inv_0
timestamp 1617951155
transform -1 0 1394 0 -1 -425
box -26 -50 13 23
use Inv  Inv_1
timestamp 1617951155
transform -1 0 1615 0 -1 -425
box -26 -50 13 23
use Inv  Inv_2
timestamp 1617951155
transform -1 0 1827 0 -1 -425
box -26 -50 13 23
use Inv  Inv_3
timestamp 1617951155
transform -1 0 2049 0 -1 -425
box -26 -50 13 23
<< labels >>
rlabel space 1014 1813 2076 1816 1 gnd
rlabel space 1014 1702 2076 1708 1 vdd
rlabel space 1014 1591 2076 1597 1 gnd
rlabel space 1014 1480 2076 1486 1 vdd
rlabel space 1014 1369 2076 1375 1 gnd
rlabel space 1014 1258 2076 1264 1 vdd
rlabel space 1014 1147 2076 1153 1 gnd
rlabel space 1014 1036 2076 1042 1 vdd
rlabel space 1014 928 2076 931 1 gnd
rlabel space 1244 66 2302 69 1 gnd
rlabel space 1244 -45 2302 -39 1 vdd
rlabel space 1244 -156 2302 -150 1 gnd
rlabel space 1244 -267 2302 -261 1 vdd
rlabel space 1244 -375 2302 -372 1 gnd
rlabel metal1 920 969 1019 973 1 Da1
rlabel metal1 1272 969 1302 973 1 Da2
rlabel metal2 1272 969 1275 1055 1 Da2
rlabel metal3 990 1052 1275 1055 1 Da2
rlabel space 920 1052 990 1055 1 Da2
rlabel metal1 1561 969 1592 973 1 Da3
rlabel metal2 1561 969 1564 1254 1 Da3
rlabel metal1 1498 1251 1564 1254 1 Da3
rlabel metal2 1413 1251 1498 1254 1 Da3
rlabel metal1 1370 1251 1413 1254 1 Da3
rlabel metal2 1347 1251 1370 1254 1 Da3
rlabel metal2 1313 1249 1317 1257 1 Da3
rlabel metal2 1313 1254 1350 1257 1 Da3
rlabel metal1 1210 1249 1317 1252 1 Da3
rlabel metal2 1122 1249 1210 1252 1 Da3
rlabel metal1 1088 1249 1122 1252 1 Da3
rlabel metal2 1064 1249 1088 1252 1 Da3
rlabel metal2 1030 1242 1033 1257 1 Da3
rlabel metal2 1030 1254 1067 1257 1 Da3
rlabel metal2 1064 1249 1067 1257 1 Da3
rlabel metal1 920 1242 1033 1245 1 Da3
rlabel metal1 1853 969 1889 973 1 Da4
rlabel metal2 1853 969 1857 1362 1 Da4
rlabel metal1 1703 1358 1857 1362 1 Da4
rlabel metal2 1552 1359 1703 1362 1 Da4
rlabel metal1 1419 1360 1552 1363 1 Da4
rlabel metal2 1252 1361 1419 1364 1 Da4
rlabel metal1 1143 1361 1252 1364 1 Da4
rlabel metal2 995 1361 1143 1364 1 Da4
rlabel metal1 920 1361 995 1364 1 Da4
rlabel metal1 975 1413 1019 1417 1 Db1
rlabel metal1 975 1413 981 1844 1 Db1
rlabel metal1 1264 1413 1302 1417 1 Db2
rlabel metal2 1264 1413 1268 1821 1 Db2
rlabel metal1 1263 1821 1267 1843 1 Db2
rlabel metal1 1554 1413 1592 1417 1 Db3
rlabel metal2 1554 1413 1558 1826 1 Db3
rlabel metal1 1554 1826 1558 1843 1 Db3
rlabel metal1 1854 1412 1889 1417 1 Db4
rlabel metal2 1854 1412 1858 1828 1 Db4
rlabel metal1 1854 1828 1858 1843 1 Db4
rlabel metal2 1017 916 1020 942 1 A1
rlabel metal2 1017 939 1219 942 1 A1
rlabel metal2 1216 939 1219 1201 1 A1
rlabel metal2 1206 1198 1219 1201 1 A1
rlabel metal2 1026 916 1029 935 1 B1
rlabel metal2 1026 932 1228 935 1 B1
rlabel metal2 1225 932 1228 1645 1 B1
rlabel metal2 1206 1642 1228 1645 1 B1
rlabel metal2 1300 916 1303 941 1 A2
rlabel metal2 1300 938 1502 941 1 A2
rlabel metal2 1498 938 1502 1201 1 A2
rlabel metal2 1489 1198 1502 1201 1 A2
rlabel metal2 1309 916 1312 934 1 B2
rlabel metal2 1309 931 1513 934 1 B2
rlabel metal2 1510 931 1513 1645 1 B2
rlabel metal2 1489 1642 1513 1645 1 B2
rlabel metal2 1592 916 1595 942 1 A3
rlabel metal2 1592 939 1790 942 1 A3
rlabel metal2 1787 939 1790 1201 1 A3
rlabel metal2 1779 1198 1790 1201 1 A3
rlabel metal2 1600 916 1603 935 1 B3
rlabel metal2 1600 932 1798 935 1 B3
rlabel metal2 1795 932 1798 1645 1 B3
rlabel metal2 1779 1642 1798 1645 1 B3
rlabel metal2 1887 914 1890 942 1 A4
rlabel metal2 1887 939 2088 942 1 A4
rlabel metal2 2085 939 2088 1201 1 A4
rlabel metal2 2076 1198 2088 1201 1 A4
rlabel metal2 1895 914 1898 934 1 B4
rlabel metal2 1895 931 2096 934 1 B4
rlabel metal2 2093 931 2096 1645 1 B4
rlabel metal2 2076 1642 2096 1645 1 B4
rlabel metal2 1118 689 1231 692 1 C0
rlabel metal1 1118 257 1122 692 1 C0
rlabel metal1 1118 257 1259 260 1 C0
rlabel metal1 1256 231 1259 260 1 C0
rlabel space 1256 209 1259 231 1 C0
rlabel space 1133 680 1228 683 1 P1
rlabel space 1134 680 1137 777 1 P1
rlabel metal2 1134 774 1213 777 1 P1
rlabel metal2 1210 774 1213 779 1 P1
rlabel metal1 1134 264 1137 683 1 P1
rlabel metal1 1134 264 1248 267 1 P1
rlabel metal2 1245 209 1248 267 1 P1
rlabel space 1126 634 1228 637 1 G1
rlabel metal1 1127 634 1130 781 1 G1
rlabel metal1 1127 778 1303 781 1 G1
rlabel m2contact 1300 778 1303 782 1 G1
rlabel space 1150 554 1228 557 1 P2
rlabel space 1150 554 1153 770 1 P2
rlabel metal2 1150 767 1496 770 1 P2
rlabel metal2 1493 767 1496 777 1 P2
rlabel metal1 1150 271 1153 557 1 P2
rlabel metal1 1150 271 1449 274 1 P2
rlabel metal2 1445 209 1448 271 1 P2
rlabel space 1141 517 1228 520 1 G2
rlabel metal1 1141 517 1144 773 1 G2
rlabel metal1 1141 770 1593 773 1 G2
rlabel metal2 1589 770 1592 780 1 G2
rlabel space 1158 404 1228 407 1 G3
rlabel metal1 1158 404 1161 766 1 G3
rlabel metal1 1158 763 1885 766 1 G3
rlabel metal2 1882 763 1885 783 1 G3
rlabel space 1166 458 1227 461 1 P3
rlabel space 1167 458 1170 763 1 P3
rlabel metal2 1167 760 1787 763 1 P3
rlabel metal2 1784 760 1787 780 1 P3
rlabel metal1 1167 277 1170 458 1 P3
rlabel metal1 1167 277 1647 280 1 P3
rlabel metal2 1644 209 1647 278 1 P3
rlabel metal3 1174 302 1195 305 1 G4
rlabel space 1174 302 1177 759 1 G4
rlabel metal1 1174 756 2181 759 1 G4
rlabel metal2 2178 756 2181 782 1 G4
rlabel metal1 1180 332 1195 335 1 P4
rlabel space 1180 332 1183 756 1 P4
rlabel metal2 1180 753 2082 756 1 P4
rlabel metal2 2079 753 2082 778 1 P4
rlabel metal1 1181 283 1184 332 1 P4
rlabel metal1 1181 283 1844 286 1 P4
rlabel metal2 1841 209 1844 283 1 P4
rlabel metal1 2043 679 2095 683 1 C1
rlabel metal1 2091 257 2095 683 1 C1
rlabel metal1 1453 257 2095 260 1 C1
rlabel space 1453 213 1456 258 1 C1
rlabel space 2043 561 2106 566 1 C2
rlabel metal1 2101 249 2105 566 1 C2
rlabel metal1 1653 249 2105 252 1 C2
rlabel space 1653 209 1656 252 1 C2
rlabel space 2043 457 2115 461 1 C3
rlabel metal1 2111 241 2115 461 1 C3
rlabel metal1 1851 241 2115 244 1 C3
rlabel space 1851 209 1854 244 1 C3
rlabel space 2062 339 2124 343 1 C4
rlabel metal1 2120 84 2124 343 1 C4
rlabel metal1 2115 84 2124 87 1 C4
rlabel space 2115 28 2118 84 1 C4
rlabel space 1894 28 1897 85 1 S4
rlabel metal2 1894 82 2038 85 1 S4
rlabel metal2 2035 82 2038 87 1 S4
rlabel space 1677 28 1680 85 1 S3
rlabel metal2 1677 82 1840 85 1 S3
rlabel metal2 1837 82 1840 87 1 S3
rlabel space 1468 28 1471 85 1 S2
rlabel metal2 1468 82 1640 85 1 S2
rlabel metal2 1637 82 1640 87 1 S2
rlabel space 1249 28 1252 85 1 S1
rlabel metal2 1249 82 1443 85 1 S1
rlabel metal2 1440 82 1443 87 1 S1
rlabel metal2 1443 -386 1447 -201 1 S1_out
rlabel metal2 1436 -204 1447 -201 1 S1_out
rlabel metal2 1660 -387 1664 -201 1 S2_out
rlabel metal2 1655 -204 1664 -201 1 S2_out
rlabel metal2 1868 -386 1872 -201 1 S3_out
rlabel metal2 1864 -204 1872 -201 1 S3_out
rlabel metal2 2085 -387 2089 -201 1 S4_out
rlabel metal2 2081 -204 2089 -201 1 S4_out
rlabel space 2313 -388 2317 -201 7 C4_out
rlabel metal2 2302 -204 2317 -201 1 C4_out
rlabel metal1 2075 -404 2089 -400 1 S4_out
rlabel metal1 2020 -404 2036 -400 1 S4_inv
rlabel metal1 1853 -404 1872 -400 1 S3_out
rlabel metal1 1800 -404 1814 -400 1 S3_inv
rlabel metal1 1641 -404 1664 -400 1 S2_out
rlabel metal1 1583 -404 1602 -400 1 S2_inv
rlabel metal1 1420 -404 1447 -400 1 S1_out
rlabel metal1 1368 -404 1381 -400 1 S1_inv
<< end >>
